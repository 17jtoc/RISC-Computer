-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Sun Feb 23 19:07:10 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY div_block IS 
	PORT
	(
		dividend :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		divisor :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		quot :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		remain :  OUT  STD_LOGIC_VECTOR(32 DOWNTO 0)
	);
END div_block;

ARCHITECTURE bdf_type OF div_block IS 

COMPONENT nonrestoring_div
	PORT(M : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 Q : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 quotient : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 remainder : OUT STD_LOGIC_VECTOR(32 DOWNTO 0)
	);
END COMPONENT;



BEGIN 



b2v_inst : nonrestoring_div
PORT MAP(M => divisor,
		 Q => dividend,
		 quotient => quot,
		 remainder => remain);


END bdf_type;